module main

import foo

println('Hello, Webpack + V.js + HMR!')
foo.hot()
