module foo

pub fn greet(msg string) {
	println('[module foo] Hello, $msg')
}
