module foo

pub fn greet(msg string) {
	println('[FOO] Hello $msg!')
}
